library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

use work.dot_fonts.all;

entity IS31FL3730_ctrl is
	port (sclk:		in std_logic;
	      kick_cmd:		in std_logic;
	      i2c_addr:		in natural;
	      module_sel:	in std_logic;
	      dot_matrix:	in dot_matrix_t;
	      device_busy:	in std_logic;

	      dbg_ps:		out natural;

	      reset_n:		out std_logic;
	      ena:		out std_logic;
	      addr:		out std_logic_vector(6 downto 0);
	      rw:		out std_logic;
	      txdata:		out std_logic_vector(7 downto 0);
	      ack_error:	buffer std_logic);
	end IS31FL3730_ctrl;

architecture arch of IS31FL3730_ctrl is
	type display_update_state is (st_ready, st_init_data_tx, st_byte_0, st_byte_1, st_byte_2, st_byte_3, st_byte_4, st_byte_5,
					st_byte_6, st_byte_7, st_end_data_tx, st_init_update, st_update_latch, st_finish);

attribute keep    :  string;
attribute mark_debug  :  string;
attribute dont_touch  :  string;

signal ns, ps		: display_update_state;

-- local signals required to latch input values when kicked
signal active_i2c_addr:	natural;
signal active_module:	std_logic;
signal active_symbol:	dot_matrix_t;

signal end_data_cnt: natural;
signal finish_cnt: natural;

attribute mark_debug of ns : signal is "TRUE";
attribute mark_debug of ps : signal is "TRUE";
attribute mark_debug of active_i2c_addr : signal is "TRUE";
attribute mark_debug of active_module : signal is "TRUE";
attribute mark_debug of active_symbol : signal is "TRUE";

attribute keep of ns : signal is "TRUE";
attribute keep of ps : signal is "TRUE";
attribute keep of active_i2c_addr : signal is "TRUE";
attribute keep of active_module : signal is "TRUE";
attribute keep of active_symbol : signal is "TRUE";

attribute dont_touch of ns : signal is "TRUE";
attribute dont_touch of ps : signal is "TRUE";
attribute dont_touch of active_i2c_addr : signal is "TRUE";
attribute dont_touch of active_module : signal is "TRUE";
attribute dont_touch of active_symbol : signal is "TRUE";


begin
	delay: process(sclk, ps)
	begin
		if rising_edge(sclk) then
			if ps = st_end_data_tx then
				end_data_cnt <= end_data_cnt + 1;
			else
				end_data_cnt <= 0;
			end if;
		end if;
	end process delay;

	sync_proc: process(sclk)
	begin
		if rising_edge(sclk) then
			-- only advance the state if the i2c controller is idle
			if device_busy = '0' or ns = st_init_data_tx or ns = st_ready then
				ps <= ns;
			end if;
			dbg_ps <= natural(display_update_state'POS(ps));
		end if;
	end process sync_proc;

	comb_proc: process(sclk, ps, kick_cmd, device_busy,
			   dot_matrix, i2c_addr, module_sel,
			   active_i2c_addr, active_module, active_symbol)
	begin
	if rising_edge(sclk) then
		case ps is
			when st_ready =>
				reset_n		<= '0';
				ena		<= '0';
				if kick_cmd = '1' then
					ns		<= st_init_data_tx; -- FIXME: make function for advancing the state ?
					active_symbol	<= dot_matrix;
					active_i2c_addr	<= i2c_addr;
					active_module 	<= module_sel;
				end if;
			when st_init_data_tx =>
				reset_n		<= '1';
				ena		<= '1';
				rw		<= '0';
				addr		<= std_logic_vector(to_unsigned(active_i2c_addr, 7));
				if active_module = '0' then
					txdata <= "00000001"; -- 0x1 mat 1 data reg address
				else
					txdata <= "00001110"; -- 0xE mat 2 data reg address
				end if;

				if device_busy = '1' then
					ns <= st_byte_0;
				end if;
			when st_byte_0 =>
				txdata		<= get_char_line(active_symbol, 0, active_module);
				if device_busy = '1' then
					ns <= st_byte_1;
				end if;
			when st_byte_1 =>
				txdata		<= get_char_line(active_symbol, 1, active_module);
				if device_busy = '1' then
					ns <= st_byte_2;
				end if;
			when st_byte_2 =>
				txdata		<= get_char_line(active_symbol, 2, active_module);
				if device_busy = '1' then
					ns <= st_byte_3;
				end if;
			when st_byte_3 =>
				txdata		<= get_char_line(active_symbol, 3, active_module);
				if device_busy = '1' then
					ns <= st_byte_4;
				end if;
			when st_byte_4 =>
				txdata		<= get_char_line(active_symbol, 4, active_module);
				if device_busy = '1' then
					ns <= st_byte_5;
				end if;
			when st_byte_5 =>
				txdata		<= get_char_line(active_symbol, 5, active_module);
				if device_busy = '1' then
					ns <= st_byte_6;
				end if;
			when st_byte_6 =>
				txdata		<= get_char_line(active_symbol, 6, active_module);
				if device_busy = '1' then
					ns <= st_byte_7;
				end if;
			when st_byte_7 =>
				txdata		<= get_char_line(active_symbol, 7, active_module);
				if device_busy = '1' then
					ns <= st_end_data_tx;
				end if;
			when st_end_data_tx =>
				ena		<= '0';
				if end_data_cnt > 200 then
					ns <= st_init_update;
				end if;
			when st_init_update =>
				ena		<= '1';
				txdata <= "00001100"; -- 0xC update reg address
				if device_busy = '1' then
					ns <= st_update_latch;
				end if;
			when st_update_latch =>
				txdata <= "11111111";
				if device_busy = '1' then
					ns <= st_finish;
				end if;
			when st_finish =>
				if finish_cnt > 200 then
					ns <= st_init_update;
				end if;
				ns <= st_ready;
		end case;
	end if;
	end process comb_proc;

end arch;
