library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

package dot_fonts is
	subtype dot_col_t is std_logic_vector(7 downto 0);

	type dot_char_t is 
		array (4 downto 0) of dot_col_t;

	function get_dot_char(ascii_code : integer) return dot_char_t;
end package dot_fonts;



package body dot_fonts is
	function get_dot_char(ascii_code : integer) return dot_char_t is
		variable dot_char : dot_char_t;
	begin
	case ascii_code is
		when 32   => dot_char := (16#00#, 16#00#, 16#00#, 16#00#, 16#00#); -- (space)
		when 33   => dot_char := (16#00#, 16#00#, 16#5f#, 16#00#, 16#00#); -- !
		when 34   => dot_char := (16#00#, 16#07#, 16#00#, 16#07#, 16#00#); -- "
		when 35   => dot_char := (16#14#, 16#7f#, 16#14#, 16#7f#, 16#14#); -- -- 
		when 36   => dot_char := (16#24#, 16#2a#, 16#7f#, 16#2a#, 16#12#); -- $
		when 37   => dot_char := (16#23#, 16#13#, 16#08#, 16#64#, 16#62#); -- %
		when 38   => dot_char := (16#36#, 16#49#, 16#55#, 16#22#, 16#50#); -- &
		when 39   => dot_char := (16#00#, 16#05#, 16#03#, 16#00#, 16#00#); -- '
		when 40   => dot_char := (16#00#, 16#1c#, 16#22#, 16#41#, 16#00#); -- (
		when 41   => dot_char := (16#00#, 16#41#, 16#22#, 16#1c#, 16#00#); -- )
		when 42   => dot_char := (16#08#, 16#2a#, 16#1c#, 16#2a#, 16#08#); -- *
		when 43   => dot_char := (16#08#, 16#08#, 16#3e#, 16#08#, 16#08#); -- +
		when 44   => dot_char := (16#00#, 16#50#, 16#30#, 16#00#, 16#00#); -- ,
		when 45   => dot_char := (16#08#, 16#08#, 16#08#, 16#08#, 16#08#); -- -
		when 46   => dot_char := (16#00#, 16#60#, 16#60#, 16#00#, 16#00#); -- .
		when 47   => dot_char := (16#20#, 16#10#, 16#08#, 16#04#, 16#02#); -- /
		when 48   => dot_char := (16#3e#, 16#51#, 16#49#, 16#45#, 16#3e#); -- 0
		when 49   => dot_char := (16#00#, 16#42#, 16#7f#, 16#40#, 16#00#); -- 1
		when 50   => dot_char := (16#42#, 16#61#, 16#51#, 16#49#, 16#46#); -- 2
		when 51   => dot_char := (16#21#, 16#41#, 16#45#, 16#4b#, 16#31#); -- 3
		when 52   => dot_char := (16#18#, 16#14#, 16#12#, 16#7f#, 16#10#); -- 4
		when 53   => dot_char := (16#27#, 16#45#, 16#45#, 16#45#, 16#39#); -- 5
		when 54   => dot_char := (16#3c#, 16#4a#, 16#49#, 16#49#, 16#30#); -- 6
		when 55   => dot_char := (16#01#, 16#71#, 16#09#, 16#05#, 16#03#); -- 7
		when 56   => dot_char := (16#36#, 16#49#, 16#49#, 16#49#, 16#36#); -- 8
		when 57   => dot_char := (16#06#, 16#49#, 16#49#, 16#29#, 16#1e#); -- 9
		when 58   => dot_char := (16#00#, 16#36#, 16#36#, 16#00#, 16#00#); -- :
		when 59   => dot_char := (16#00#, 16#56#, 16#36#, 16#00#, 16#00#); -- ;
		when 60   => dot_char := (16#00#, 16#08#, 16#14#, 16#22#, 16#41#); -- <
		when 61   => dot_char := (16#14#, 16#14#, 16#14#, 16#14#, 16#14#); -- =
		when 62   => dot_char := (16#41#, 16#22#, 16#14#, 16#08#, 16#00#); -- >
		when 63   => dot_char := (16#02#, 16#01#, 16#51#, 16#09#, 16#06#); -- ?
		when 64   => dot_char := (16#32#, 16#49#, 16#79#, 16#41#, 16#3e#); -- @
		when 65   => dot_char := (16#7e#, 16#11#, 16#11#, 16#11#, 16#7e#); -- A
		when 66   => dot_char := (16#7f#, 16#49#, 16#49#, 16#49#, 16#36#); -- B
		when 67   => dot_char := (16#3e#, 16#41#, 16#41#, 16#41#, 16#22#); -- C
		when 68   => dot_char := (16#7f#, 16#41#, 16#41#, 16#22#, 16#1c#); -- D
		when 69   => dot_char := (16#7f#, 16#49#, 16#49#, 16#49#, 16#41#); -- E
		when 70   => dot_char := (16#7f#, 16#09#, 16#09#, 16#01#, 16#01#); -- F
		when 71   => dot_char := (16#3e#, 16#41#, 16#41#, 16#51#, 16#32#); -- G
		when 72   => dot_char := (16#7f#, 16#08#, 16#08#, 16#08#, 16#7f#); -- H
		when 73   => dot_char := (16#00#, 16#41#, 16#7f#, 16#41#, 16#00#); -- I
		when 74   => dot_char := (16#20#, 16#40#, 16#41#, 16#3f#, 16#01#); -- J
		when 75   => dot_char := (16#7f#, 16#08#, 16#14#, 16#22#, 16#41#); -- K
		when 76   => dot_char := (16#7f#, 16#40#, 16#40#, 16#40#, 16#40#); -- L
		when 77   => dot_char := (16#7f#, 16#02#, 16#04#, 16#02#, 16#7f#); -- M
		when 78   => dot_char := (16#7f#, 16#04#, 16#08#, 16#10#, 16#7f#); -- N
		when 79   => dot_char := (16#3e#, 16#41#, 16#41#, 16#41#, 16#3e#); -- O
		when 80   => dot_char := (16#7f#, 16#09#, 16#09#, 16#09#, 16#06#); -- P
		when 81   => dot_char := (16#3e#, 16#41#, 16#51#, 16#21#, 16#5e#); -- Q
		when 82   => dot_char := (16#7f#, 16#09#, 16#19#, 16#29#, 16#46#); -- R
		when 83   => dot_char := (16#46#, 16#49#, 16#49#, 16#49#, 16#31#); -- S
		when 84   => dot_char := (16#01#, 16#01#, 16#7f#, 16#01#, 16#01#); -- T
		when 85   => dot_char := (16#3f#, 16#40#, 16#40#, 16#40#, 16#3f#); -- U
		when 86   => dot_char := (16#1f#, 16#20#, 16#40#, 16#20#, 16#1f#); -- V
		when 87   => dot_char := (16#7f#, 16#20#, 16#18#, 16#20#, 16#7f#); -- W
		when 88   => dot_char := (16#63#, 16#14#, 16#08#, 16#14#, 16#63#); -- X
		when 89   => dot_char := (16#03#, 16#04#, 16#78#, 16#04#, 16#03#); -- Y
		when 90   => dot_char := (16#61#, 16#51#, 16#49#, 16#45#, 16#43#); -- Z
		when 91   => dot_char := (16#00#, 16#00#, 16#7f#, 16#41#, 16#41#); -- (
		when 92   => dot_char := (16#02#, 16#04#, 16#08#, 16#10#, 16#20#); -- \
		when 93   => dot_char := (16#41#, 16#41#, 16#7f#, 16#00#, 16#00#); -- )
		when 94   => dot_char := (16#04#, 16#02#, 16#01#, 16#02#, 16#04#); -- ^
		when 95   => dot_char := (16#40#, 16#40#, 16#40#, 16#40#, 16#40#); -- _
		when 96   => dot_char := (16#00#, 16#01#, 16#02#, 16#04#, 16#00#); -- `
		when 97   => dot_char := (16#20#, 16#54#, 16#54#, 16#54#, 16#78#); -- a
		when 98   => dot_char := (16#7f#, 16#48#, 16#44#, 16#44#, 16#38#); -- b
		when 99   => dot_char := (16#38#, 16#44#, 16#44#, 16#44#, 16#20#); -- c
		when 100  => dot_char := (16#38#, 16#44#, 16#44#, 16#48#, 16#7f#); -- d
		when 101  => dot_char := (16#38#, 16#54#, 16#54#, 16#54#, 16#18#); -- e
		when 102  => dot_char := (16#08#, 16#7e#, 16#09#, 16#01#, 16#02#); -- f
		when 103  => dot_char := (16#08#, 16#14#, 16#54#, 16#54#, 16#3c#); -- g
		when 104  => dot_char := (16#7f#, 16#08#, 16#04#, 16#04#, 16#78#); -- h
		when 105  => dot_char := (16#00#, 16#44#, 16#7d#, 16#40#, 16#00#); -- i
		when 106  => dot_char := (16#20#, 16#40#, 16#44#, 16#3d#, 16#00#); -- j
		when 107  => dot_char := (16#00#, 16#7f#, 16#10#, 16#28#, 16#44#); -- k
		when 108  => dot_char := (16#00#, 16#41#, 16#7f#, 16#40#, 16#00#); -- l
		when 109  => dot_char := (16#7c#, 16#04#, 16#18#, 16#04#, 16#78#); -- m
		when 110  => dot_char := (16#7c#, 16#08#, 16#04#, 16#04#, 16#78#); -- n
		when 111  => dot_char := (16#38#, 16#44#, 16#44#, 16#44#, 16#38#); -- o
		when 112  => dot_char := (16#7c#, 16#14#, 16#14#, 16#14#, 16#08#); -- p
		when 113  => dot_char := (16#08#, 16#14#, 16#14#, 16#18#, 16#7c#); -- q
		when 114  => dot_char := (16#7c#, 16#08#, 16#04#, 16#04#, 16#08#); -- r
		when 115  => dot_char := (16#48#, 16#54#, 16#54#, 16#54#, 16#20#); -- s
		when 116  => dot_char := (16#04#, 16#3f#, 16#44#, 16#40#, 16#20#); -- t
		when 117  => dot_char := (16#3c#, 16#40#, 16#40#, 16#20#, 16#7c#); -- u
		when 118  => dot_char := (16#1c#, 16#20#, 16#40#, 16#20#, 16#1c#); -- v
		when 119  => dot_char := (16#3c#, 16#40#, 16#30#, 16#40#, 16#3c#); -- w
		when 120  => dot_char := (16#44#, 16#28#, 16#10#, 16#28#, 16#44#); -- x
		when 121  => dot_char := (16#0c#, 16#50#, 16#50#, 16#50#, 16#3c#); -- y
		when 122  => dot_char := (16#44#, 16#64#, 16#54#, 16#4c#, 16#44#); -- z
		when 123  => dot_char := (16#00#, 16#08#, 16#36#, 16#41#, 16#00#); -- {
		when 124  => dot_char := (16#00#, 16#00#, 16#7f#, 16#00#, 16#00#); -- |
		when 125  => dot_char := (16#00#, 16#41#, 16#36#, 16#08#, 16#00#); -- }
		when 126  => dot_char := (16#08#, 16#08#, 16#2a#, 16#1c#, 16#08#); -- ~
		when others => dot_char := (16#ff#, 16#ff#, 16#ff#, 16#ff#, 16#ff#); -- (undefined)
	end case;
	return dot_char;
	end function get_dot_char;

end package body dot_fonts;
